library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control is
    port(
        clk: in std_logic; --sygnał zegarowy
        reset : in std_logic; 
        IR: in signed(15 downto 0);
        Salu : out signed(4 downto 0);
        S_ALU_A, S_ALU_B, S_ALU_Y: out signed(3 downto 0); -- sygnały sterujące [Salu] [SBB] [SBC] [SBA]
        Sid, Sadr: out signed(2 downto 0);
        Smar, Smbr, WR, RD: out std_logic
    );
end entity;

architecture rtl of control is
    type state_type is (fetch, fetch2, decode, mov, mov2, mov3, add, add2, add3, add4, add5,
    sub, sub2, sub3, sub4, sub5, cmpA, cmpA_2, cmpA_3, cmpA_4, cmpR, push, pop, pop2, pop3, oxnorR, oxnorC,
    rpl8A, rpl8A_2, rpl8A_3, rpl8A_4, rpl8A_5, rpl8R, rpl4A, rpl4A_2, rpl4A_3, rpl4A_4, rpl4A_5, rpl4R );
    signal state : state_type;

    begin
    process (clk, reset)
        begin
            if(reset = '1') then
                state <= fetch;
            elsif (clk'event and clk = '1') then
                case state is
                    when fetch =>
                        state <= fetch2;
                    when fetch2 =>
                        state <= decode;
                    --dekodowanie rozkazu procesora
                    when decode =>
                        -- pierwsze 2 bity - ilość argumentów operacji
                        case IR(15 downto 14) is
                            -- jednoargumentowe
                            when "01" =>
                                case IR(13 downto 11) is
                                    when "000" =>
                                        state <= push;
                                    when "001" =>
                                        state <= pop;
                                    when "010" =>
                                        if IR(10) = '0' then
                                            state <= rpl8A;
                                        else
                                            state <= rpl8R;
                                        end if;
                                    when "011" =>
                                        if IR(10) = '0' then
                                            state <= rpl4A;
                                        else
                                            state <= rpl4R;
                                        end if;
                                    when others =>
                                        state <= fetch;
                                end case;
                            --dwuargumentowe: arg1 - adres, arg2 - rejestr lub arg1 - rejestr, arg2 - rejestr
                            when "10" =>
                                case IR(13 downto 11) is
                                    when "000" =>
                                        state <= mov;
                                    when "001" =>
                                        state <= add;
                                    when "010" =>
                                        state <= sub;
                                    when "011" =>
                                        if (IR(10) = '0') then
                                            state <= cmpA;
                                        else 
                                            state <= cmpR;
                                        end if;
                                    when "100" =>
                                        if (IR(10) = '0') then
                                            state <= oxnorC;
                                        else 
                                            state <= oxnorR;
                                        end if;
                                    when others =>
                                        state <= fetch;
                                end case;
                            when others =>
                                state <= fetch;
                        end case;
                    when push =>
                        state <= fetch;
                    when pop =>
                        state <= pop2;
                    when pop2 =>
                        state <= pop3;
                    when pop3 =>
                        state <= fetch;
                    when rpl8A =>
                        state <= rpl8A_2;
                    when rpl8A_2 =>
                        state <= rpl8A_3;
                    when rpl8A_3 =>
                        state <= rpl8A_4;
                    when rpl8A_4 =>
                        state <= rpl8A_5;
                    when rpl8A_5 =>
                        state <= fetch;
                    when rpl8R =>
                        state <= fetch;
                    when rpl4A =>
                        state <= rpl4A_2;
                    when rpl4A_2 =>
                        state <= rpl4A_3;
                    when rpl4A_3 =>
                        state <= rpl4A_4;
                    when rpl4A_4 =>
                        state <= rpl4A_5;
                    when rpl4A_5 =>
                        state <= fetch;
                    when rpl4R =>
                        state <= fetch;
                    when mov =>
                        state <= mov2;
                    when mov2 => 
                        state <= mov3;
                    when mov3 =>
                        state <= fetch;
                    when add =>
                        state <= add2;
                    when add2 =>
                        state <= add3;
                    when add3 =>
                        state <= add4;
                    when add4 =>
                        state <= add5;
                    when add5 =>
                        state <= fetch;
                    when sub =>
                        state <= sub2;
                    when sub2 =>
                        state <= sub3;
                    when sub3 =>
                        state <= sub4;
                    when sub4 =>
                        state <= sub5;
                    when sub5 =>
                        state <= fetch;
                    when cmpA =>
                        state <= cmpA_2;
                    when cmpA_2 =>
                        state <= cmpA_3;
                    when cmpA_3 =>
                        state <= cmpA_4;
                    when cmpA_4 =>
                        state <= fetch;
                    when cmpR =>
                        state <= fetch;
                    when oxnorC =>
                        state <= fetch;
                    when oxnorR =>
                        state <= fetch;
                    when others =>
                        state <= fetch;
                end case;
            end if;
    end process;

    process(state)
    begin
        case state is
            when fetch => --wystaw zawartość rejestru PC -> ADR -> MAR
                Sadr <= "001";                  -- PC -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              -- nic nie rób (tu było psute)
                Sid <= "001";                   -- PC++
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR  
                WR <= '0';                      -- nie zapisuj do RAM 
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when fetch2 => --odczytaj zawartość komórki pamięci RAM spod adresu wskazywanego przez MAR i umieść ją w MBR, MBR -> DATA_INPUT -> ALU_A -> ALU_Y -> IR
                Sadr <= "000";                  -- AD -> ADR            - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= "0000";              -- ALU_Y -> IR
                Sid <= "000";                   -- nic nie rób
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when decode => --dekodowanie rozkazu przechowywanego w rejestrze IR
                Sadr <= "000";                  -- AD -> ADR            - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A  - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B  - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              -- nie rób nic          
                Sid <= "000";                   -- nie rób nic          
                Smar <= '0';                    -- pamiętanie MAR       
                Smbr <= '0';                    -- pamiętanie MBR       
                WR <= '0';                      -- nie zapisuj do RAM   
                RD <= '0';                      -- nie odczytuj z RAM   
                Salu <= "00000";                -- ALU_A -> ALU_Y       - nie ma znaczenia co tutaj będzie
            when push => --dodawanie wartości na stos (do RAMu pod adres wskazany przez rejetr SP), dekrementacja SP, 
                Sadr <= "010";                  -- SP -> ADR
                S_ALU_A <= IR(3 downto 0);      -- REG(X) -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              -- nie zapisuj ALU_Y do rejestru
                Sid <= "011";                   -- SP--
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '1';                    -- ALU_Y -> MBR
                WR <= '1';                      -- zapisz zawartość MBR do RAM
                RD <= '0';                      -- nie odczytuj z RAM
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when pop => --zwiększ wskaźnik stosu o 1
                Sadr <= "000";                  -- AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              -- nic nie rób
                Sid <= "010";                   -- SP++
                Smar <= '0';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '0';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when pop2 => --ustaw rejestr MAR na wartość spod wskaźnika szczytu stosu zwiększonego o 1
                Sadr <= "010";                  -- AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              -- nic nie rób
                Sid <= "000";                   -- nic nie rób
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y            - nie ma znaczenia co tutaj będzie
            when pop3 => --odczytaj wartosc na szczycie stosu w pamięci RAM i wprowadź odczytaną wartość do rejestru
                Sadr <= "000";                  -- AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= IR(3 downto 0);      -- ALU_Y -> REJ
                Sid <= "000";                   -- nic nie rób
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y  
            when rpl8A => --pierwsza część pobierania adresu z pamięci - wystawienie zawartości PC na ADR
                Sadr <= "001";                  -- PC -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              -- pamiętanie ALU_Y      -bez znaczenia
                Sid <= "001";                   -- PC++
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y  
            when rpl8A_2 => --wprowadzenie odczytanej wartości do rejestru rozkazów IR
                Sadr <= "000";                  -- AD -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B   -bez znaczenia
                S_ALU_Y <= "0000";              -- ALU_Y -> IR
                Sid <= "000";                   -- nic nie rób
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when rpl8A_3 => --wystawienie zawartości IR na ADR, a następnie na MAR
                Sadr <= "100";                  -- IR -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              -- nie rób nic
                Sid <= "000";                   -- nie rób nic
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y
            when rpl8A_4 => --odczytanie zawartości RAM spod adresu umieszczonego w MAR oraz obliczenie wyniku operacji
                Sadr <= "000";                  -- AD -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B   -bez znaczenia
                S_ALU_Y <= "1111";              -- nie zapisuj do rejestru
                Sid <= "000";                   -- nie rób nic
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "10110";                -- RPL8(ALU_A) -> ALU_Y
            when rpl8A_5 => --zapisanie obliczonego wyniku operacji do pamięci RAM
                Sadr <= "000";                  -- AD -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_Y <= "1111";              -- nie zapisuj do rejestru
                Sid <= "000";                   -- nie rób nic
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '1';                    -- ALU_Y -> MBR
                WR <= '1';                      -- zapisz zawartość MBR do RAM
                RD <= '0';                      -- nie odczytuj z RAM
                Salu <= "11111";                -- nie rób nic
            when rpl8R => --odczytanie podanego w rozkazie rejestru i przesłanie jego zawartości do wejścia ALU_A, wykonanie operacji RPL8, przesłanie wyniku operacji do rejestru 
                Sadr <= "000";                  -- AD -> ADR
                S_ALU_A <= IR(3 downto 0);      -- REJ -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= IR(3 downto 0);      -- ALU_Y -> REJ
                Sid <= "000";                   --nie rób nic
                Smar <= '0';                    -- pamiętanie MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '0';                      -- nie odczytuj z RAM
                Salu <= "10110";                -- RPL8(ALU_A) -> ALU_Y
            when rpl4A => --pierwsza część pobierania adresu z pamięci - wystawienie zawartości PC na ADR
                Sadr <= "001";                  -- PC -> ADR
                S_ALU_A <= "0000";              -- DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              -- DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              -- pamiętanie ALU_Y      -bez znaczenia
                Sid <= "001";                   -- PC++
                Smar <= '1';                    -- ADR -> MAR
                Smbr <= '0';                    -- pamiętanie MBR
                WR <= '0';                      -- nie zapisuj do RAM
                RD <= '1';                      -- RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                -- ALU_A -> ALU_Y  
            when rpl4A_2 => --wprowadzenie odczytanej wartości do rejestru rozkazów IR
                Sadr <= "000";                  --AD -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   -bez znaczenia
                S_ALU_Y <= "0000";              --ALU_Y -> IR
                Sid <= "000";                   --nic nie rób
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when rpl4A_3 => --wystawienie zawartości IR na ADR, a następnie na MAR
                Sadr <= "100";                  --IR -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              --nie rób nic
                Sid <= "000";                   --nie rób nic
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when rpl4A_4 => --odczytanie zawartości RAM spod adresu umieszczonego w MAR oraz obliczenie wyniku operacji
                Sadr <= "000";                  --AD -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   -bez znaczenia
                S_ALU_Y <= "1111";              --nie zapisuj do rejestru
                Sid <= "000";                   --nie rób nic
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "10111";                --RPL4(ALU_A) -> ALU_Y
            when rpl4A_5 => --zapisanie obliczonego wyniku operacji do pamięci RAM
                Sadr <= "000";                  --AD -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_Y <= "1111";              --nie zapisuj do rejestru
                Sid <= "000";                   --nie rób nic
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '1';                    --ALU_Y -> MBR
                WR <= '1';                      --zapisz zawartość MBR do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "11111";                --nie rób nic
            when rpl4R => --odczytanie podanego w rozkazie rejestru i przesłanie jego zawartości do wejścia ALU_A, wykonanie operacji RPL4, przesłanie wyniku operacji do rejestru 
                Sadr <= "000";                  --AD -> ADR
                S_ALU_A <= IR(3 downto 0);      --REJ -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B
                S_ALU_Y <= IR(3 downto 0);      --ALU_Y -> REJ
                Sid <= "000";                   --nie rób nic
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "10111";                --RPL4(ALU_A) -> ALU_Y
            when mov => --zapis zawartości rejestru do TMP, pierwsza część pobierania adresu z pamięci (czyli argumentu operacji mov)
                Sadr <= "001";                  --PC -> ADR
                S_ALU_A <= IR(3 downto 0);      --REJ -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie 
                S_ALU_Y <= "0001";              --ALU_Y -> TMP
                Sid <= "001";                   --zwiększ PC o 1
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --Nie zapisuj do RAM 
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when mov2 => --wprowadzenie pobranego adresu z pamięci do rejestru rozkazów IR
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "0000";              --ALU_Y -> IR
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when mov3 => --zapisanie zawartości TMP do komórki pamięci RAM o adresie podanym w IR
                Sadr <= "100";                  --IR -> ADR
                S_ALU_A <= "0001";              --TMP -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '1';                    --ALU_Y -> MBR
                WR <= '1';                      --zapisz zawartość MBR do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "00000";                --ALU_A -> ALU_Y            - nie ma znaczenia co tutaj będzie
            when add => --zapis zawartości rejestru do TMP, pierwsza część pobierania adresu z pamięci (czyli argumentu operacji add)
                Sadr <= "001";                  --PC -> ADR
                S_ALU_A <= IR(3 downto 0);      --REJ -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie      
                S_ALU_Y <= "0001";              --ALU_Y -> TMP
                Sid <= "001";                   --zwiększ PC o 1
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --Nie zapisuj do RAM 
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when add2 => --wprowadzenie pobranego adresu z pamięci do rejestru rozkazów IR
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "0000";              --ALU_Y -> IR
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when add3 => --pobieranie zawartości komórki RAM spod adresu będącego argumentem operacji 
                Sadr <= "100";                  --IR -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y            - nie ma znaczenia co tutaj będzie
            when add4 => --dodanie obu wartości do siebie
                Sadr <= "000";                  --AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0001";              --TMP -> ALU_B
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00010";                --ALU_A + ALU_B -> ALU_Y
            when add5 => --zapisanie wyniku z ALU_Y do MBR, a następnie do RAM
                Sadr <= "000";                  --AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '1';                    --ALU_Y -> MBR
                WR <= '1';                      --zapisz zawartość MBR do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "11111";                --pamiętanie zawartości ALU_Y
            when sub => --zapis zawartości rejestru do TMP, pierwsza część pobierania adresu z pamięci (czyli argumentu operacji sub)
                Sadr <= "001";                  --PC -> ADR
                S_ALU_A <= IR(3 downto 0);      --REJ -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie      
                S_ALU_Y <= "0001";              --ALU_Y -> TMP
                Sid <= "001";                   --zwiększ PC o 1
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --Nie zapisuj do RAM 
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when sub2 => --wprowadzenie pobranego adresu z pamięci do rejestru rozkazów IR
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "0000";              --ALU_Y -> IR
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when sub3 => --pobieranie zawartości komórki RAM spod adresu będącego argumentem operacji
                Sadr <= "100";                  --IR -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y            - nie ma znaczenia co tutaj będzie
            when sub4 => --odjęcie obu wartości od siebie
                Sadr <= "000";                  --AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0001";              --TMP -> ALU_B
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00011";                --ALU_A - ALU_B -> ALU_Y
            when sub5 => --zapisanie wyniku z ALU_Y do MBR, a następnie do RAM
                Sadr <= "000";                  --AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '1';                    --ALU_Y -> MBR
                WR <= '1';                      --zapisz zawartość MBR do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "11111";                --pamiętanie zawartości ALU_Y
            when cmpA => --zapis zawartości rejestru do TMP, pierwsza część pobierania adresu z pamięci (czyli argumentu operacji cmp)
                Sadr <= "001";                  --PC -> ADR
                S_ALU_A <= IR(3 downto 0);      --REJ -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie      
                S_ALU_Y <= "0001";              --ALU_Y -> TMP
                Sid <= "001";                   --zwiększ PC o 1
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --Nie zapisuj do RAM 
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when cmpA_2 => --wprowadzenie pobranego adresu z pamięci do rejestru rozkazów IR
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B   - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "0000";              --ALU_Y -> IR
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y
            when cmpA_3 => --pobieranie zawartości komórki RAM spod adresu będącego argumentem operacji 
                Sadr <= "100";                  --IR -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A       - nie ma znaczenia co tutaj będzie
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B       - nie ma znaczenia co tutaj będzie
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '1';                    --ADR -> MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "00000";                --ALU_A -> ALU_Y            - nie ma znaczenia co tutaj będzie
            when cmpA_4 => --porównanie wartości i ustawienie flag ALU
                Sadr <= "000";                  --AD -> ADR                 - nie ma znaczenia co tutaj będzie
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0001";              --TMP -> ALU_B
                S_ALU_Y <= "1111";              --nie zapisuj ALU_Y do rejestru
                Sid <= "000";                   --nic nie zmieniaj w PC, SP i AD
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '1';                      --RAM -> MBR -> DATA_INPUT
                Salu <= "10101";                --CMP(ALU_A, ALU_B) -> ALU_Y
            when cmpR =>  --pobranie wartości ze wskazanych rejestrów (REJ1 -> ALU_A, REJ2 -> ALU_B), porównanie wartości, ustawienie flag ALU
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= IR(7 downto 4);      --REJ1 -> ALU_A
                S_ALU_B <= IR(3 downto 0);      --REJ2 -> ALU_B
                S_ALU_Y <= "1111";              --nic nie rób
                Sid <= "000";                   --nic nie rób
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "10101";                --CMP(ALU_A, ALU_B) -> ALU_Y
            when oxnorC => --obliczenie xnor dla rejestru i stałej oraz zapisanie wyniku do rejestru (REJ1 -> ALU_A, )
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tu będzie
                S_ALU_A <= IR(8 downto 5);      --REJ1 -> ALU_A
                S_ALU_B <= "1010";              --STAŁA -> ALU_B
                S_ALU_Y <= IR(8 downto 5);      --ALU_Y -> REJ1
                Sid <= "000";                   --nic nie rób
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "00111";                --XNOR(REJ1, STAŁA) -> ALU_Y
            when oxnorR => --obliczenie xnor dla dwóch rejestrów oraz zapisanie wyniku do pierwszego z rejestów (REJ1 -> ALU_A, REJ2 -> ALU_B, ALU_Y -> REJ1)
                Sadr <= "000";                  --AD -> ADR             - nie ma znaczenia co tutaj będzie
                S_ALU_A <= IR(7 downto 4);      --REJ1 -> ALU_A
                S_ALU_B <= IR(3 downto 0);      --REJ2 -> ALU_B
                S_ALU_Y <= IR(7 downto 4);      --ALU_Y -> REJ1
                Sid <= "000";                   --nic nie rób
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "00111";                --XNOR(REJ1, REJ2) -> ALU_Y
            when others => --gdy nie rozpoznano rozkazu
                Sadr <= "000";                  --AD -> ADR
                S_ALU_A <= "0000";              --DATA_INPUT -> ALU_A
                S_ALU_B <= "0000";              --DATA_INPUT -> ALU_B
                S_ALU_Y <= "1111";              --nic nie rób
                Sid <= "000";                   --nic nie rób
                Smar <= '0';                    --pamiętanie MAR
                Smbr <= '0';                    --pamiętanie MBR
                WR <= '0';                      --nie zapisuj do RAM
                RD <= '0';                      --nie odczytuj z RAM
                Salu <= "11111";                --pamiętanie ALU_Y      - nie ma znaczenia co tutaj będzie
        end case;
    end process;
end rtl;